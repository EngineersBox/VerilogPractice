module q2_fsm #(parameter BIT_WIDTH = 32)(bitstring);
	input [BIT_WIDTH - 1 : 0] bitstring;



endmodule
